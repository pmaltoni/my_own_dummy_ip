pmaltoni@lagrev3.ee.ethz.ch.42609:1599369532